netcdf partition_metadata_3 {
dimensions:
	NX = 6 ;
	NY = 4 ;
	P = 3 ;
	L = 2 ;
	R = 2 ;
	B = UNLIMITED ; // (0 currently)
	T = UNLIMITED ; // (0 currently)

group: bounding_boxes {
  variables:
  	int domain_x(P) ;
  	int domain_extent_x(P) ;
  	int domain_y(P) ;
  	int domain_extent_y(P) ;
  data:

   domain_x = 0, 2, 4 ;

   domain_extent_x = 2, 2, 2 ;

   domain_y = 0, 0, 0 ;

   domain_extent_y = 4, 4, 4 ;
  } // group bounding_boxes

group: connectivity {
  variables:
  	int left_neighbours(P) ;
  	int left_neighbour_ids(L) ;
  	int left_neighbour_halos(L) ;
  	int right_neighbours(P) ;
  	int right_neighbour_ids(R) ;
  	int right_neighbour_halos(R) ;
  	int bottom_neighbours(P) ;
  	int bottom_neighbour_ids(B) ;
  	int bottom_neighbour_halos(B) ;
  	int top_neighbours(P) ;
  	int top_neighbour_ids(T) ;
  	int top_neighbour_halos(T) ;
  data:

   left_neighbours = 0, 1, 1 ;

   left_neighbour_ids = 0, 1 ;

   left_neighbour_halos = 4, 4 ;

   right_neighbours = 1, 1, 0 ;

   right_neighbour_ids = 1, 2 ;

   right_neighbour_halos = 4, 4 ;

   bottom_neighbours = 0, 0, 0 ;

   top_neighbours = 0, 0, 0 ;
  } // group connectivity
}
