netcdf rect3030.res {

group: structure {

  // group attributes:
  		:type = "simple_rectangular" ;
  } // group structure

group: data {
  dimensions:
  	x = 30 ;
  	y = 30 ;
  	nLayers = 1 ;
  variables:
  	double mask(x, y) ;
  	double cice(x, y) ;
  		cice:missing_value = -2.03703597633449e+90 ;
  	double hice(x, y) ;
  		hice:missing_value = -2.03703597633449e+90 ;
  	double hsnow(x, y) ;
  		hsnow:missing_value = -2.03703597633449e+90 ;
  	double sss(x, y) ;
  		sss:missing_value = -2.03703597633449e+90 ;
  	double sst(x, y) ;
  		sst:missing_value = -2.03703597633449e+90 ;
  	double tice(x, y, nLayers) ;
  		tice:missing_value = -2.03703597633449e+90 ;
  data:

   mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      0, 0, 0, 0, 0, 0,
  0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      0, 0, 0, 0, 0, 0,
  0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 
      0, 0, 0, 0, 0, 0,
  0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 
      0, 0, 0, 0, 0, 0,
  0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      1, 0, 0, 0, 0, 0,
  1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      1, 1, 0, 0, 0, 0,
  0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      1, 0, 0, 0, 0, 0,
  0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      1, 1, 0, 0, 0, 0,
  0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 
      0, 1, 1, 0, 0, 0,
  1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 
      1, 1, 0, 0, 0, 0,
  1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 
      1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      1, 1, 0, 0, 0, 0,
  1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      1, 1, 0, 0, 0, 0,
  1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
      1, 0, 0, 0, 0, 0,
  1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 
      1, 0, 0, 0, 0, 0,
  1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 
      1, 0, 0, 0, 0, 0,
  1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 
      0, 0, 0, 0, 0, 0 ;

   cice =
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.1, 0, 0, 0, 0, 0, 0.1, 
      0.1, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0.1, 0.1, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.1, 0.1, 0.2, 0.2, 0.1, 0.1, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0.1, 0.1, 0.2, 0.3, 
      0.4, 0.5, 0.4, 0.3, 0.3, 0.2, 0.2, 0.3, 0.2, 0.1, 0.1, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0.1, 0.2, 0.4, 0.5, 0.6, 0.5, 0.5, 0.4, 
      0.3, 0.3, 0.4, 0.2, 0.1, 0.1, -2.03703597633449e+90, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, 0.1, 0.2, 0.5, 0.7, 
      0.8, 0.7, 0.8, 0.6, 0.4, 0.5, 0.3, 0.2, 0.2, 0.1, 0.1, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.3, 0.5, 0.7, 0.9, 0.9, 0.9, 0.8, 0.6, 0.8, 0.6, 0.4, 0.2, 0.1, 0.1, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.6, 
      -2.03703597633449e+90, 0.7, 0.8, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.8, 
      0.5, 0.3, 0.2, 0.1, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.6, -2.03703597633449e+90, 0.8, 0.8, 0.9, 0.9, 
      0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.7, 0.5, 0.4, 0.2, 0.1, 0.1, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.7, 0.8, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 
      0.9, 0.9, 0.6, 0.5, 0.3, 0.2, 0.1, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.8, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.6, 0.5, 
      0.3, 0.1, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.9, -2.03703597633449e+90, 0.8, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 
      0.9, 0.9, 0.9, 0.8, -2.03703597633449e+90, 0.4, 0.3, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.9, 0.9, 0.9, 0.8, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.7, 0.5, 0.3, 0.1, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.8, 0.9, 0.9, 0.9, 0.7, 0.6, 0.4, 0.3, 0.2, 0.1, 0.1, 0.1, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, 0, 0.9, 0.9, 0.9, 0.9, 0.9, 0.8, 
      0.7, 0.5, 0.3, 0.2, 0.2, 0.1, 0.1, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.9, 0.7, 0.5, 0.3, 0.3, 0.4, 0.2, 0.1, 0.1, 0, 
      0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.6, 0.5, 0.5, 0.4, 0.3, 0.2, 0.2, 0.2, 0.1, 0, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.4, 0.2, 0.1, 0.1, 0.2, 0.1, 0.1, 0.1, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.3, 0.2, 0.1, -2.03703597633449e+90, 0.1, 0, 0, 0, 0, 
      -2.03703597633449e+90, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.2, 0.1, 0, 0, -2.03703597633449e+90, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.3, 0.2, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.2, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.2, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90 ;

   hice =
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.2, 0, 0, 0, 0, 0, 0.2, 
      0.2, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.2, 0.2, 0.2, 0.2, 0.2, 
      0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0.2, 0.2, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.2, 0.2, 0.4, 0.4, 0.2, 0.2, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0.2, 0.2, 0.4, 0.6, 
      0.8, 1, 0.8, 0.6, 0.6, 0.4, 0.4, 0.6, 0.4, 0.2, 0.2, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0.2, 0.4, 0.8, 1, 1.2, 1, 1, 0.8, 0.6, 
      0.6, 0.8, 0.4, 0.2, 0.2, -2.03703597633449e+90, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, 0.2, 0.4, 1, 1.4, 1.6, 
      1.4, 1.6, 1.2, 0.8, 1, 0.6, 0.4, 0.4, 0.2, 0.2, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.6, 1, 1.4, 1.8, 1.8, 1.8, 1.6, 1.2, 1.6, 1.2, 0.8, 0.4, 0.2, 0.2, 0, 
      0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 1.2, 
      -2.03703597633449e+90, 1.4, 1.6, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.6, 1, 
      0.6, 0.4, 0.2, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 1.2, -2.03703597633449e+90, 1.6, 1.6, 1.8, 1.8, 
      1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.4, 1, 0.8, 0.4, 0.2, 0.2, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, 1.4, 1.6, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 
      1.8, 1.8, 1.2, 1, 0.6, 0.4, 0.2, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      1.6, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.2, 1, 
      0.6, 0.2, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      1.8, -2.03703597633449e+90, 1.6, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 
      1.8, 1.8, 1.8, 1.6, -2.03703597633449e+90, 0.8, 0.6, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      1.8, 1.8, 1.8, 1.6, 1.8, 1.8, 1.8, 1.8, 1.8, 1.8, 1.4, 1, 0.6, 0.2, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      1.6, 1.8, 1.8, 1.8, 1.4, 1.2, 0.8, 0.6, 0.4, 0.2, 0.2, 0.2, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, 0, 1.8, 1.8, 1.8, 1.8, 1.8, 1.6, 
      1.4, 1, 0.6, 0.4, 0.4, 0.2, 0.2, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 1.8, 1.4, 1, 0.6, 0.6, 0.8, 0.4, 0.2, 0.2, 0, 0, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 1.2, 1, 1, 0.8, 0.6, 0.4, 0.4, 0.4, 0.2, 0, 0, 
      0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.8, 0.4, 0.2, 0.2, 0.4, 0.2, 0.2, 0.2, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.6, 0.4, 0.2, -2.03703597633449e+90, 0.2, 0, 0, 0, 0, 
      -2.03703597633449e+90, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.4, 0.2, 0, 0, -2.03703597633449e+90, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.6, 0.4, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.4, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.4, 0.2, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90 ;

   hsnow =
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.05, 0, 0, 0, 0, 0, 
      0.05, 0.05, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.05, 0.05, 0.05, 0.05, 
      0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0.05, 0.05, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.05, 0.05, 0.1, 0.1, 0.05, 
      0.05, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0.05, 0.05, 0.1, 0.15, 
      0.2, 0.25, 0.2, 0.15, 0.15, 0.1, 0.1, 0.15, 0.1, 0.05, 0.05, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0.05, 0.1, 0.2, 0.25, 0.3, 0.25, 0.25, 
      0.2, 0.15, 0.15, 0.2, 0.1, 0.05, 0.05, -2.03703597633449e+90, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, 0.05, 0.1, 0.25, 0.35, 
      0.4, 0.35, 0.4, 0.3, 0.2, 0.25, 0.15, 0.1, 0.1, 0.05, 0.05, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.15, 0.25, 0.35, 0.45, 0.45, 0.45, 0.4, 0.3, 0.4, 0.3, 0.2, 0.1, 0.05, 
      0.05, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0.3, 
      -2.03703597633449e+90, 0.35, 0.4, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 
      0.4, 0.25, 0.15, 0.1, 0.05, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.3, -2.03703597633449e+90, 0.4, 0.4, 0.45, 
      0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.35, 0.25, 0.2, 0.1, 0.05, 
      0.05, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.35, 0.4, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 
      0.45, 0.45, 0.45, 0.3, 0.25, 0.15, 0.1, 0.05, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.4, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 
      0.3, 0.25, 0.15, 0.05, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.45, -2.03703597633449e+90, 0.4, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 
      0.45, 0.45, 0.45, 0.45, 0.4, -2.03703597633449e+90, 0.2, 0.15, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.45, 0.45, 0.45, 0.4, 0.45, 0.45, 0.45, 0.45, 0.45, 0.45, 0.35, 0.25, 
      0.15, 0.05, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.4, 0.45, 0.45, 0.45, 0.35, 0.3, 0.2, 0.15, 0.1, 0.05, 0.05, 0.05, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, 0, 0.45, 0.45, 0.45, 0.45, 0.45, 
      0.4, 0.35, 0.25, 0.15, 0.1, 0.1, 0.05, 0.05, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.45, 0.35, 0.25, 0.15, 0.15, 0.2, 0.1, 0.05, 
      0.05, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.3, 0.25, 0.25, 0.2, 0.15, 0.1, 0.1, 0.1, 0.05, 
      0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.2, 0.1, 0.05, 0.05, 0.1, 0.05, 0.05, 0.05, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.15, 0.1, 0.05, -2.03703597633449e+90, 0.05, 0, 0, 0, 0, 
      -2.03703597633449e+90, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.1, 0.05, 0, 0, -2.03703597633449e+90, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.15, 0.1, 0.05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0.1, 0.05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.1, 0.05, 0.05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0.05, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90 ;

   sss =
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 
      32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 
      32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, -2.03703597633449e+90, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, -2.03703597633449e+90, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 32, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, -2.03703597633449e+90, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      32, -2.03703597633449e+90, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 32, 
      32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  32, -2.03703597633449e+90, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, -2.03703597633449e+90, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  32, 32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, -2.03703597633449e+90, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  32, 32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  32, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  32, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, -2.03703597633449e+90, -2.03703597633449e+90, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  32, -2.03703597633449e+90, -2.03703597633449e+90, 32, 32, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  32, 32, 32, 32, 32, 32, 32, 32, -2.03703597633449e+90, 32, 32, 32, 32, 
      32, 32, 32, 32, 32, 32, -2.03703597633449e+90, -2.03703597633449e+90, 
      32, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90 ;

   sst =
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -0.2, 0, 0, 0, 0, 0, 
      -0.2, -0.2, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -0.2, -0.2, -0.2, -0.2, 
      -0.2, -0.2, -0.2, -0.2, -0.2, -0.2, -0.2, -0.2, -0.2, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -0.2, -0.2, -0.4, -0.4, -0.4, -0.4, -0.4, -0.4, -0.2, -0.2, -0.4, -0.4, 
      -0.2, -0.2, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, -0.2, -0.2, -0.4, 
      -0.6, -0.8, -1, -0.8, -0.6, -0.6, -0.4, -0.4, -0.6, -0.4, -0.2, -0.2, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, -0.2, -0.4, -0.8, -1, -1.2, -1, -1, -0.8, 
      -0.6, -0.6, -0.8, -0.4, -0.2, -0.2, -2.03703597633449e+90, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -0.2, -0.4, -1, -1.4, 
      -1.6, -1.4, -1.6, -1.2, -0.8, -1, -0.6, -0.4, -0.4, -0.2, -0.2, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -0.6, -1, -1.4, -1.8, -1.8, -1.8, -1.6, -1.2, -1.6, -1.2, -0.8, -0.4, 
      -0.2, -0.2, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -1.2, 
      -2.03703597633449e+90, -1.4, -1.6, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, 
      -1.6, -1, -0.6, -0.4, -0.2, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -1.2, -2.03703597633449e+90, -1.6, -1.6, -1.8, 
      -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.4, -1, -0.8, -0.4, -0.2, 
      -0.2, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -1.4, -1.6, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, 
      -1.8, -1.8, -1.8, -1.2, -1, -0.6, -0.4, -0.2, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -1.6, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, 
      -1.2, -1, -0.6, -0.2, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -1.8, -2.03703597633449e+90, -1.6, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, 
      -1.8, -1.8, -1.8, -1.8, -1.6, -2.03703597633449e+90, -0.8, -0.6, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -1.8, -1.8, -1.8, -1.6, -1.8, -1.8, -1.8, -1.8, -1.8, -1.8, -1.4, -1, 
      -0.6, -0.2, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -1.6, -1.8, -1.8, -1.8, -1.4, -1.2, -0.8, -0.6, -0.4, -0.2, -0.2, -0.2, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, 0, 0, 0, 0, -1.8, -1.8, -1.8, -1.8, -1.8, 
      -1.6, -1.4, -1, -0.6, -0.4, -0.4, -0.2, -0.2, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -1.8, -1.4, -1, -0.6, -0.6, -0.8, -0.4, -0.2, 
      -0.2, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -1.2, -1, -1, -0.8, -0.6, -0.4, -0.4, -0.4, 
      -0.2, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -0.8, -0.4, -0.2, -0.2, -0.4, -0.2, -0.2, -0.2, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -0.6, -0.4, -0.2, -2.03703597633449e+90, -0.2, 0, 0, 0, 0, 
      -2.03703597633449e+90, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -0.4, -0.2, 0, 0, -2.03703597633449e+90, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -0.6, -0.4, -0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -0.4, -0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -0.4, -0.2, -0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -0.2, 0, 0, 0, 0, 0, 0, 0, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90,
  0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90,
  0, 0, 0, 0, 0, 0, 0, 0, -2.03703597633449e+90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, -2.03703597633449e+90, -2.03703597633449e+90, 0, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90, -2.03703597633449e+90, 
      -2.03703597633449e+90, -2.03703597633449e+90 ;

   tice =
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.6,
  -0.6,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -0.6,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.6,
  -0.6,
  -0.7,
  -0.7,
  -0.7,
  -0.7,
  -0.7,
  -0.7,
  -0.6,
  -0.6,
  -0.7,
  -0.7,
  -0.6,
  -0.6,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.6,
  -0.6,
  -0.7,
  -0.8,
  -0.9,
  -1,
  -0.9,
  -0.8,
  -0.8,
  -0.7,
  -0.7,
  -0.8,
  -0.7,
  -0.6,
  -0.6,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.6,
  -0.7,
  -0.9,
  -1,
  -1.1,
  -1,
  -1,
  -0.9,
  -0.8,
  -0.8,
  -0.9,
  -0.7,
  -0.6,
  -0.6,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -0.6,
  -0.7,
  -1,
  -1.2,
  -1.3,
  -1.2,
  -1.3,
  -1.1,
  -0.9,
  -1,
  -0.8,
  -0.7,
  -0.7,
  -0.6,
  -0.6,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.8,
  -1,
  -1.2,
  -1.4,
  -1.4,
  -1.4,
  -1.3,
  -1.1,
  -1.3,
  -1.1,
  -0.9,
  -0.7,
  -0.6,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.1,
  -2.03703597633449e+90,
  -1.2,
  -1.3,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.3,
  -1,
  -0.8,
  -0.7,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.1,
  -2.03703597633449e+90,
  -1.3,
  -1.3,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.2,
  -1,
  -0.9,
  -0.7,
  -0.6,
  -0.6,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.2,
  -1.3,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.1,
  -1,
  -0.8,
  -0.7,
  -0.6,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.3,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.1,
  -1,
  -0.8,
  -0.6,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.4,
  -2.03703597633449e+90,
  -1.3,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.3,
  -2.03703597633449e+90,
  -0.9,
  -0.8,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.4,
  -1.4,
  -1.4,
  -1.3,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.2,
  -1,
  -0.8,
  -0.6,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.3,
  -1.4,
  -1.4,
  -1.4,
  -1.2,
  -1.1,
  -0.9,
  -0.8,
  -0.7,
  -0.6,
  -0.6,
  -0.6,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.4,
  -1.3,
  -1.2,
  -1,
  -0.8,
  -0.7,
  -0.7,
  -0.6,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.4,
  -1.2,
  -1,
  -0.8,
  -0.8,
  -0.9,
  -0.7,
  -0.6,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -1.1,
  -1,
  -1,
  -0.9,
  -0.8,
  -0.7,
  -0.7,
  -0.7,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.9,
  -0.7,
  -0.6,
  -0.6,
  -0.7,
  -0.6,
  -0.6,
  -0.6,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.8,
  -0.7,
  -0.6,
  -2.03703597633449e+90,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.7,
  -0.6,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.8,
  -0.7,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.7,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.7,
  -0.6,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.6,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -0.5,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90,
  -2.03703597633449e+90 ;
  } // group data
}
